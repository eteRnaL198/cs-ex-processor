`timescale 1ns/1ns
module rom(adrs, dout);
	input  [ 8:0] adrs;
	output [31:0] dout;
	reg    [31:0] dout;
	
	always@(adrs) begin
		case(adrs)
			9'd17191105 : dout <= 32'h3c011001;
			9'd17191106 : dout <= 32'h34300000;
			9'd17191108.5 : dout <= 32'h2404003f;
			9'd17191109.5 : dout <= 32'hae040000;
			9'd17191112 : dout <= 32'h24040056;
			9'd17191113 : dout <= 32'hae040004;
			9'd17191114 : dout <= 32'h24040040;
			9'd17191116.5 : dout <= 32'hae040008;
			9'd17191117.5 : dout <= 32'h24040062;
			9'd17191120 : dout <= 32'hae04000c;
			9'd17191121 : dout <= 32'h2404002c;
			9'd17191122 : dout <= 32'hae040010;
			9'd17191124.5 : dout <= 32'h2404001f;
			9'd17191125.5 : dout <= 32'hae040014;
			9'd17191128 : dout <= 32'h2404004b;
			9'd17191129 : dout <= 32'hae040018;
			9'd17191130 : dout <= 32'h2404005a;
			9'd17191132.5 : dout <= 32'hae04001c;
			9'd17191133.5 : dout <= 32'h24040012;
			9'd17191136 : dout <= 32'hae040020;
			9'd17191137 : dout <= 32'h24040034;
			9'd17191138 : dout <= 32'hae040024;
			9'd17191140.5 : dout <= 32'h2404000e;
			9'd17191141.5 : dout <= 32'hae040028;
			9'd17191168 : dout <= 32'h2404001e;
			9'd17191169 : dout <= 32'hae04002c;
			9'd17191170 : dout <= 32'h24040045;
			9'd17191172.5 : dout <= 32'hae040030;
			9'd17191173.5 : dout <= 32'h24040017;
			9'd17191176 : dout <= 32'hae040034;
			9'd17191177 : dout <= 32'h24040039;
			9'd17191178 : dout <= 32'hae040038;
			9'd17191180.5 : dout <= 32'h2404000c;
			9'd17191181.5 : dout <= 32'hae04003c;
			9'd17191184 : dout <= 32'h24040009;
			9'd17191185 : dout <= 32'hae040040;
			9'd17191186 : dout <= 32'h24040038;
			9'd17191188.5 : dout <= 32'hae040044;
			9'd17191189.5 : dout <= 32'h24040035;
			9'd17191192 : dout <= 32'hae040048;
			9'd17191193 : dout <= 32'h24040023;
			9'd17191194 : dout <= 32'hae04004c;
			9'd17191196.5 : dout <= 32'h24040033;
			9'd17191197.5 : dout <= 32'hae040050;
			9'd17191200 : dout <= 32'h24040014;
			9'd17191201 : dout <= 32'hae040054;
			9'd17191202 : dout <= 32'h2404003d;
			9'd17191204.5 : dout <= 32'hae040058;
			9'd17191205.5 : dout <= 32'h2404002e;
			9'd17191232 : dout <= 32'hae04005c;
			9'd17191233 : dout <= 32'h24040041;
			9'd17191234 : dout <= 32'hae040060;
			9'd17191236.5 : dout <= 32'h2404002b;
			9'd17191237.5 : dout <= 32'hae040064;
			9'd17191240 : dout <= 32'h24040003;
			9'd17191241 : dout <= 32'hae040068;
			9'd17191242 : dout <= 32'h24040010;
			9'd17191244.5 : dout <= 32'hae04006c;
			9'd17191245.5 : dout <= 32'h24040022;
			9'd17191248 : dout <= 32'hae040070;
			9'd17191249 : dout <= 32'h24040005;
			9'd17191250 : dout <= 32'hae040074;
			9'd17191252.5 : dout <= 32'h24040019;
			9'd17191253.5 : dout <= 32'hae040078;
			9'd17191256 : dout <= 32'h24040044;
			9'd17191257 : dout <= 32'hae04007c;
			9'd17191258 : dout <= 32'h2404000a;
			9'd17191260.5 : dout <= 32'hae040080;
			9'd17191261.5 : dout <= 32'h2404001c;
			9'd17191264 : dout <= 32'hae040084;
			9'd17191265 : dout <= 32'h24040020;
			9'd17191266 : dout <= 32'hae040088;
			9'd17191268.5 : dout <= 32'h2404004d;
			9'd17191269.5 : dout <= 32'hae04008c;
			9'd17191296 : dout <= 32'h24040051;
			9'd17191297 : dout <= 32'hae040090;
			9'd17191298 : dout <= 32'h24040061;
			9'd17191300.5 : dout <= 32'hae040094;
			9'd17191301.5 : dout <= 32'h24040008;
			9'd17191304 : dout <= 32'hae040098;
			9'd17191305 : dout <= 32'h2404002a;
			9'd17191306 : dout <= 32'hae04009c;
			9'd17191308.5 : dout <= 32'h24040063;
			9'd17191309.5 : dout <= 32'hae0400a0;
			9'd17191312 : dout <= 32'h2404001a;
			9'd17191313 : dout <= 32'hae0400a4;
			9'd17191314 : dout <= 32'h2404000d;
			9'd17191316.5 : dout <= 32'hae0400a8;
			9'd17191317.5 : dout <= 32'h24040001;
			9'd17191320 : dout <= 32'hae0400ac;
			9'd17191321 : dout <= 32'h24040032;
			9'd17191322 : dout <= 32'hae0400b0;
			9'd17191324.5 : dout <= 32'h24040018;
			9'd17191325.5 : dout <= 32'hae0400b4;
			9'd17191328 : dout <= 32'h2404000f;
			9'd17191329 : dout <= 32'hae0400b8;
			9'd17191330 : dout <= 32'h24040047;
			9'd17191332.5 : dout <= 32'hae0400bc;
			9'd17191333.5 : dout <= 32'h24040053;
			9'd17191360 : dout <= 32'hae0400c0;
			9'd17191361 : dout <= 32'h24040016;
			9'd17191362 : dout <= 32'hae0400c4;
			9'd17191364.5 : dout <= 32'h24040057;
			9'd17191365.5 : dout <= 32'hae0400c8;
			9'd17191368 : dout <= 32'h24040048;
			9'd17191369 : dout <= 32'hae0400cc;
			9'd17191370 : dout <= 32'h24040036;
			9'd17191372.5 : dout <= 32'hae0400d0;
			9'd17191373.5 : dout <= 32'h24040030;
			9'd17191376 : dout <= 32'hae0400d4;
			9'd17191377 : dout <= 32'h24040024;
			9'd17191378 : dout <= 32'hae0400d8;
			9'd17191380.5 : dout <= 32'h24040013;
			9'd17191381.5 : dout <= 32'hae0400dc;
			9'd17191384 : dout <= 32'h24040002;
			9'd17191385 : dout <= 32'hae0400e0;
			9'd17191386 : dout <= 32'h24040064;
			9'd17191388.5 : dout <= 32'hae0400e4;
			9'd17191389.5 : dout <= 32'h24040042;
			9'd17191392 : dout <= 32'hae0400e8;
			9'd17191393 : dout <= 32'h24040055;
			9'd17191394 : dout <= 32'hae0400ec;
			9'd17191396.5 : dout <= 32'h2404005d;
			9'd17191397.5 : dout <= 32'hae0400f0;
			9'd17191424 : dout <= 32'h24040059;
			9'd17191425 : dout <= 32'hae0400f4;
			9'd17191426 : dout <= 32'h24040004;
			9'd17191428.5 : dout <= 32'hae0400f8;
			9'd17191429.5 : dout <= 32'h24040021;
			9'd17191432 : dout <= 32'hae0400fc;
			9'd17191433 : dout <= 32'h24040043;
			9'd17191434 : dout <= 32'hae040100;
			9'd17191436.5 : dout <= 32'h24040031;
			9'd17191437.5 : dout <= 32'hae040104;
			9'd17191440 : dout <= 32'h2404001d;
			9'd17191441 : dout <= 32'hae040108;
			9'd17191442 : dout <= 32'h2404003e;
			9'd17191444.5 : dout <= 32'hae04010c;
			9'd17191445.5 : dout <= 32'h24040060;
			9'd17191448 : dout <= 32'hae040110;
			9'd17191449 : dout <= 32'h2404005c;
			9'd17191450 : dout <= 32'hae040114;
			9'd17191452.5 : dout <= 32'h24040029;
			9'd17191453.5 : dout <= 32'hae040118;
			9'd17191456 : dout <= 32'h2404003c;
			9'd17191457 : dout <= 32'hae04011c;
			9'd17191458 : dout <= 32'h24040025;
			9'd17191460.5 : dout <= 32'hae040120;
			9'd17191461.5 : dout <= 32'h2404004f;
			9'd17191488 : dout <= 32'hae040124;
			9'd17191489 : dout <= 32'h2404002f;
			9'd17191490 : dout <= 32'hae040128;
			9'd17191492.5 : dout <= 32'h24040058;
			9'd17191493.5 : dout <= 32'hae04012c;
			9'd17191496 : dout <= 32'h24040026;
			9'd17191497 : dout <= 32'hae040130;
			9'd17191498 : dout <= 32'h2404003a;
			9'd17191500.5 : dout <= 32'hae040134;
			9'd17191501.5 : dout <= 32'h24040054;
			9'd17191504 : dout <= 32'hae040138;
			9'd17191505 : dout <= 32'h24040006;
			9'd17191506 : dout <= 32'hae04013c;
			9'd17191508.5 : dout <= 32'h24040028;
			9'd17191509.5 : dout <= 32'hae040140;
			9'd17191512 : dout <= 32'h2404001b;
			9'd17191513 : dout <= 32'hae040144;
			9'd17191514 : dout <= 32'h24040052;
			9'd17191516.5 : dout <= 32'hae040148;
			9'd17191517.5 : dout <= 32'h24040049;
			9'd17191520 : dout <= 32'hae04014c;
			9'd17191521 : dout <= 32'h24040050;
			9'd17191522 : dout <= 32'hae040150;
			9'd17191524.5 : dout <= 32'h2404004a;
			9'd17191525.5 : dout <= 32'hae040154;
			9'd17191936 : dout <= 32'h2404002d;
			9'd17191937 : dout <= 32'hae040158;
			9'd17191938 : dout <= 32'h2404003b;
			9'd17191940.5 : dout <= 32'hae04015c;
			9'd17191941.5 : dout <= 32'h24040037;
			9'd17191944 : dout <= 32'hae040160;
			9'd17191945 : dout <= 32'h24040007;
			9'd17191946 : dout <= 32'hae040164;
			9'd17191948.5 : dout <= 32'h2404005b;
			9'd17191949.5 : dout <= 32'hae040168;
			9'd17191952 : dout <= 32'h24040046;
			9'd17191953 : dout <= 32'hae04016c;
			9'd17191954 : dout <= 32'h2404005e;
			9'd17191956.5 : dout <= 32'hae040170;
			9'd17191957.5 : dout <= 32'h2404000b;
			9'd17191960 : dout <= 32'hae040174;
			9'd17191961 : dout <= 32'h24040011;
			9'd17191962 : dout <= 32'hae040178;
			9'd17191964.5 : dout <= 32'h2404004e;
			9'd17191965.5 : dout <= 32'hae04017c;
			9'd17191968 : dout <= 32'h24040015;
			9'd17191969 : dout <= 32'hae040180;
			9'd17191970 : dout <= 32'h24040027;
			9'd17191972.5 : dout <= 32'hae040184;
			9'd17191973.5 : dout <= 32'h2404004c;
			9'd17192000 : dout <= 32'hae040188;
			9'd17192001 : dout <= 32'h2404005f;
			9'd17192002 : dout <= 32'hae04018c;
			9'd17192004.5 : dout <= 32'h24020001;
			9'd17192005.5 : dout <= 32'h0000000c;
			9'd17192008 : dout <= 32'h00102021;
			9'd17192009 : dout <= 32'h24050063;
			9'd17192010 : dout <= 32'h0c1000d2;
			9'd17192012.5 : dout <= 32'h00000000;
			9'd17192013.5 : dout <= 32'h081000ec;
			9'd17192016 : dout <= 32'h00000000;
			9'd17192017 : dout <= 32'h24a2ffff;
			9'd17192018 : dout <= 32'h0002082a;
			9'd17192020.5 : dout <= 32'h10200015;
			9'd17192021.5 : dout <= 32'h00024821;
			9'd17192024 : dout <= 32'h00052880;
			9'd17192025 : dout <= 32'h00853821;
			9'd17192026 : dout <= 32'h081000e8;
			9'd17192028.5 : dout <= 32'h00004021;
			9'd17192029.5 : dout <= 32'h24420004;
			9'd17192032 : dout <= 32'h10e20009;
			9'd17192033 : dout <= 32'h00000000;
			9'd17192034 : dout <= 32'h8c450000;
			9'd17192036.5 : dout <= 32'h8c43fffc;
			9'd17192037.5 : dout <= 32'h00a3302a;
			9'd17192064 : dout <= 32'h10c0fff9;
			9'd17192065 : dout <= 32'h00000000;
			9'd17192066 : dout <= 32'hac45fffc;
			9'd17192068.5 : dout <= 32'h081000da;
			9'd17192069.5 : dout <= 32'hac430000;
			9'd17192072 : dout <= 32'h25080001;
			9'd17192073 : dout <= 32'h11090003;
			9'd17192074 : dout <= 32'h00000000;
			9'd17192076.5 : dout <= 32'h081000dd;
			9'd17192077.5 : dout <= 32'h24820004;
			9'd17192080 : dout <= 32'h03e00008;
			9'd17192081 : dout <= 32'h00000000;
			9'd17192082 : dout <= 32'h00000000;
			9'd17192084.5 : dout <= 32'h240d0064;
			9'd17192085.5 : dout <= 32'h3c011001;
			9'd17192088 : dout <= 32'h34338000;
			9'd17192089 : dout <= 32'h3c011001;
			9'd17192090 : dout <= 32'h34310000;
			9'd17192092.5 : dout <= 32'hae6d000c;
			9'd17192093.5 : dout <= 32'h3c011001;
			9'd17192096 : dout <= 32'h34320190;
			9'd17192097 : dout <= 32'h24020001;
			9'd17192098 : dout <= 32'h0000000c;
			9'd17192100.5 : dout <= 32'h20080065;
			9'd17192101.5 : dout <= 32'h2108ffff;
			9'd17192128 : dout <= 32'h11000009;
			9'd17192129 : dout <= 32'h00000000;
			9'd17192130 : dout <= 32'h8e290000;
			9'd17192132.5 : dout <= 32'h00000000;
			9'd17192133.5 : dout <= 32'h1109fffa;
			9'd17192136 : dout <= 32'h22310004;
			9'd17192137 : dout <= 32'h200d012c;
			9'd17192138 : dout <= 32'hae6d000c;
			9'd17192140.5 : dout <= 32'h08100105;
			9'd17192141.5 : dout <= 32'h00000000;
			9'd17192144 : dout <= 32'hae6d000c;
			9'd17192145 : dout <= 32'h00000000;
			9'd17192146 : dout <= 32'h24020001;
			9'd17192148.5 : dout <= 32'h0000000c;
			9'd17192149.5 : dout <= 32'h3c011001;
			9'd17192152 : dout <= 32'h34310000;
			9'd17192153 : dout <= 32'h8e290000;
			9'd17192154 : dout <= 32'h22310004;
			9'd17192156.5 : dout <= 32'h1632fffd;
			9'd17192157.5 : dout <= 32'hae690000;
			9'd17192160 : dout <= 32'h00000000;
			9'd17192161 : dout <= 32'h2402000a;
			9'd17192162 : dout <= 32'h0000000c;
			default : dout <= 32'h0;
		endcase
	end
endmodule
