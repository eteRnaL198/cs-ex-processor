`timescale 1ns/1ns
module rom(adrs, dout);
	input  [ 8:0] adrs;
	output [31:0] dout;
	reg    [31:0] dout;
	
	always@(adrs) begin
		case(adrs)
			9'd0 : dout <= 32'h3c011001;
			9'd1 : dout <= 32'h34300000;
			9'd2 : dout <= 32'h2404003f;
			9'd3 : dout <= 32'hae040000;
			9'd4 : dout <= 32'h24040056;
			9'd5 : dout <= 32'hae040004;
			9'd6 : dout <= 32'h24040040;
			9'd7 : dout <= 32'hae040008;
			9'd8 : dout <= 32'h24040062;
			9'd9 : dout <= 32'hae04000c;
			9'd10 : dout <= 32'h2404002c;
			9'd11 : dout <= 32'hae040010;
			9'd12 : dout <= 32'h2404001f;
			9'd13 : dout <= 32'hae040014;
			9'd14 : dout <= 32'h2404004b;
			9'd15 : dout <= 32'hae040018;
			9'd16 : dout <= 32'h2404005a;
			9'd17 : dout <= 32'hae04001c;
			9'd18 : dout <= 32'h24040012;
			9'd19 : dout <= 32'hae040020;
			9'd20 : dout <= 32'h24040034;
			9'd21 : dout <= 32'hae040024;
			9'd22 : dout <= 32'h2404000e;
			9'd23 : dout <= 32'hae040028;
			9'd24 : dout <= 32'h2404001e;
			9'd25 : dout <= 32'hae04002c;
			9'd26 : dout <= 32'h24040045;
			9'd27 : dout <= 32'hae040030;
			9'd28 : dout <= 32'h24040017;
			9'd29 : dout <= 32'hae040034;
			9'd30 : dout <= 32'h24040039;
			9'd31 : dout <= 32'hae040038;
			9'd32 : dout <= 32'h2404000c;
			9'd33 : dout <= 32'hae04003c;
			9'd34 : dout <= 32'h24040009;
			9'd35 : dout <= 32'hae040040;
			9'd36 : dout <= 32'h24040038;
			9'd37 : dout <= 32'hae040044;
			9'd38 : dout <= 32'h24040035;
			9'd39 : dout <= 32'hae040048;
			9'd40 : dout <= 32'h24040023;
			9'd41 : dout <= 32'hae04004c;
			9'd42 : dout <= 32'h24040033;
			9'd43 : dout <= 32'hae040050;
			9'd44 : dout <= 32'h24040014;
			9'd45 : dout <= 32'hae040054;
			9'd46 : dout <= 32'h2404003d;
			9'd47 : dout <= 32'hae040058;
			9'd48 : dout <= 32'h2404002e;
			9'd49 : dout <= 32'hae04005c;
			9'd50 : dout <= 32'h24040041;
			9'd51 : dout <= 32'hae040060;
			9'd52 : dout <= 32'h2404002b;
			9'd53 : dout <= 32'hae040064;
			9'd54 : dout <= 32'h24040003;
			9'd55 : dout <= 32'hae040068;
			9'd56 : dout <= 32'h24040010;
			9'd57 : dout <= 32'hae04006c;
			9'd58 : dout <= 32'h24040022;
			9'd59 : dout <= 32'hae040070;
			9'd60 : dout <= 32'h24040005;
			9'd61 : dout <= 32'hae040074;
			9'd62 : dout <= 32'h24040019;
			9'd63 : dout <= 32'hae040078;
			9'd64 : dout <= 32'h24040044;
			9'd65 : dout <= 32'hae04007c;
			9'd66 : dout <= 32'h2404000a;
			9'd67 : dout <= 32'hae040080;
			9'd68 : dout <= 32'h2404001c;
			9'd69 : dout <= 32'hae040084;
			9'd70 : dout <= 32'h24040020;
			9'd71 : dout <= 32'hae040088;
			9'd72 : dout <= 32'h2404004d;
			9'd73 : dout <= 32'hae04008c;
			9'd74 : dout <= 32'h24040051;
			9'd75 : dout <= 32'hae040090;
			9'd76 : dout <= 32'h24040061;
			9'd77 : dout <= 32'hae040094;
			9'd78 : dout <= 32'h24040008;
			9'd79 : dout <= 32'hae040098;
			9'd80 : dout <= 32'h2404002a;
			9'd81 : dout <= 32'hae04009c;
			9'd82 : dout <= 32'h24040063;
			9'd83 : dout <= 32'hae0400a0;
			9'd84 : dout <= 32'h2404001a;
			9'd85 : dout <= 32'hae0400a4;
			9'd86 : dout <= 32'h2404000d;
			9'd87 : dout <= 32'hae0400a8;
			9'd88 : dout <= 32'h24040001;
			9'd89 : dout <= 32'hae0400ac;
			9'd90 : dout <= 32'h24040032;
			9'd91 : dout <= 32'hae0400b0;
			9'd92 : dout <= 32'h24040018;
			9'd93 : dout <= 32'hae0400b4;
			9'd94 : dout <= 32'h2404000f;
			9'd95 : dout <= 32'hae0400b8;
			9'd96 : dout <= 32'h24040047;
			9'd97 : dout <= 32'hae0400bc;
			9'd98 : dout <= 32'h24040053;
			9'd99 : dout <= 32'hae0400c0;
			9'd100 : dout <= 32'h24040016;
			9'd101 : dout <= 32'hae0400c4;
			9'd102 : dout <= 32'h24040057;
			9'd103 : dout <= 32'hae0400c8;
			9'd104 : dout <= 32'h24040048;
			9'd105 : dout <= 32'hae0400cc;
			9'd106 : dout <= 32'h24040036;
			9'd107 : dout <= 32'hae0400d0;
			9'd108 : dout <= 32'h24040030;
			9'd109 : dout <= 32'hae0400d4;
			9'd110 : dout <= 32'h24040024;
			9'd111 : dout <= 32'hae0400d8;
			9'd112 : dout <= 32'h24040013;
			9'd113 : dout <= 32'hae0400dc;
			9'd114 : dout <= 32'h24040002;
			9'd115 : dout <= 32'hae0400e0;
			9'd116 : dout <= 32'h24040064;
			9'd117 : dout <= 32'hae0400e4;
			9'd118 : dout <= 32'h24040042;
			9'd119 : dout <= 32'hae0400e8;
			9'd120 : dout <= 32'h24040055;
			9'd121 : dout <= 32'hae0400ec;
			9'd122 : dout <= 32'h2404005d;
			9'd123 : dout <= 32'hae0400f0;
			9'd124 : dout <= 32'h24040059;
			9'd125 : dout <= 32'hae0400f4;
			9'd126 : dout <= 32'h24040004;
			9'd127 : dout <= 32'hae0400f8;
			9'd128 : dout <= 32'h24040021;
			9'd129 : dout <= 32'hae0400fc;
			9'd130 : dout <= 32'h24040043;
			9'd131 : dout <= 32'hae040100;
			9'd132 : dout <= 32'h24040031;
			9'd133 : dout <= 32'hae040104;
			9'd134 : dout <= 32'h2404001d;
			9'd135 : dout <= 32'hae040108;
			9'd136 : dout <= 32'h2404003e;
			9'd137 : dout <= 32'hae04010c;
			9'd138 : dout <= 32'h24040060;
			9'd139 : dout <= 32'hae040110;
			9'd140 : dout <= 32'h2404005c;
			9'd141 : dout <= 32'hae040114;
			9'd142 : dout <= 32'h24040029;
			9'd143 : dout <= 32'hae040118;
			9'd144 : dout <= 32'h2404003c;
			9'd145 : dout <= 32'hae04011c;
			9'd146 : dout <= 32'h24040025;
			9'd147 : dout <= 32'hae040120;
			9'd148 : dout <= 32'h2404004f;
			9'd149 : dout <= 32'hae040124;
			9'd150 : dout <= 32'h2404002f;
			9'd151 : dout <= 32'hae040128;
			9'd152 : dout <= 32'h24040058;
			9'd153 : dout <= 32'hae04012c;
			9'd154 : dout <= 32'h24040026;
			9'd155 : dout <= 32'hae040130;
			9'd156 : dout <= 32'h2404003a;
			9'd157 : dout <= 32'hae040134;
			9'd158 : dout <= 32'h24040054;
			9'd159 : dout <= 32'hae040138;
			9'd160 : dout <= 32'h24040006;
			9'd161 : dout <= 32'hae04013c;
			9'd162 : dout <= 32'h24040028;
			9'd163 : dout <= 32'hae040140;
			9'd164 : dout <= 32'h2404001b;
			9'd165 : dout <= 32'hae040144;
			9'd166 : dout <= 32'h24040052;
			9'd167 : dout <= 32'hae040148;
			9'd168 : dout <= 32'h24040049;
			9'd169 : dout <= 32'hae04014c;
			9'd170 : dout <= 32'h24040050;
			9'd171 : dout <= 32'hae040150;
			9'd172 : dout <= 32'h2404004a;
			9'd173 : dout <= 32'hae040154;
			9'd174 : dout <= 32'h2404002d;
			9'd175 : dout <= 32'hae040158;
			9'd176 : dout <= 32'h2404003b;
			9'd177 : dout <= 32'hae04015c;
			9'd178 : dout <= 32'h24040037;
			9'd179 : dout <= 32'hae040160;
			9'd180 : dout <= 32'h24040007;
			9'd181 : dout <= 32'hae040164;
			9'd182 : dout <= 32'h2404005b;
			9'd183 : dout <= 32'hae040168;
			9'd184 : dout <= 32'h24040046;
			9'd185 : dout <= 32'hae04016c;
			9'd186 : dout <= 32'h2404005e;
			9'd187 : dout <= 32'hae040170;
			9'd188 : dout <= 32'h2404000b;
			9'd189 : dout <= 32'hae040174;
			9'd190 : dout <= 32'h24040011;
			9'd191 : dout <= 32'hae040178;
			9'd192 : dout <= 32'h2404004e;
			9'd193 : dout <= 32'hae04017c;
			9'd194 : dout <= 32'h24040015;
			9'd195 : dout <= 32'hae040180;
			9'd196 : dout <= 32'h24040027;
			9'd197 : dout <= 32'hae040184;
			9'd198 : dout <= 32'h2404004c;
			9'd199 : dout <= 32'hae040188;
			9'd200 : dout <= 32'h2404005f;
			9'd201 : dout <= 32'hae04018c;
			9'd202 : dout <= 32'h24020001;
			9'd203 : dout <= 32'h0000000c;
			9'd204 : dout <= 32'h00102021;
			9'd205 : dout <= 32'h24050063;
			9'd206 : dout <= 32'h0c1000d2;
			9'd207 : dout <= 32'h00000000;
			9'd208 : dout <= 32'h081000da;
			9'd209 : dout <= 32'h00000000;
			9'd210 : dout <= 32'h00001021;
			9'd211 : dout <= 32'hac800000;
			9'd212 : dout <= 32'h24420001;
			9'd213 : dout <= 32'h00a2182a;
			9'd214 : dout <= 32'h1060fffc;
			9'd215 : dout <= 32'h24840004;
			9'd216 : dout <= 32'h03e00008;
			9'd217 : dout <= 32'h00000000;
			9'd218 : dout <= 32'h00000000;
			9'd219 : dout <= 32'h240d0064;
			9'd220 : dout <= 32'h3c011001;
			9'd221 : dout <= 32'h34338000;
			9'd222 : dout <= 32'h3c011001;
			9'd223 : dout <= 32'h34310000;
			9'd224 : dout <= 32'hae6d000c;
			9'd225 : dout <= 32'h3c011001;
			9'd226 : dout <= 32'h34320190;
			9'd227 : dout <= 32'h24020001;
			9'd228 : dout <= 32'h0000000c;
			9'd229 : dout <= 32'h20080065;
			9'd230 : dout <= 32'h2108ffff;
			9'd231 : dout <= 32'h11000009;
			9'd232 : dout <= 32'h00000000;
			9'd233 : dout <= 32'h8e290000;
			9'd234 : dout <= 32'h00000000;
			9'd235 : dout <= 32'h1109fffa;
			9'd236 : dout <= 32'h22310004;
			9'd237 : dout <= 32'h200d012c;
			9'd238 : dout <= 32'hae6d000c;
			9'd239 : dout <= 32'h081000f3;
			9'd240 : dout <= 32'h00000000;
			9'd241 : dout <= 32'hae6d000c;
			9'd242 : dout <= 32'h00000000;
			9'd243 : dout <= 32'h24020001;
			9'd244 : dout <= 32'h0000000c;
			9'd245 : dout <= 32'h3c011001;
			9'd246 : dout <= 32'h34310000;
			9'd247 : dout <= 32'h8e290000;
			9'd248 : dout <= 32'h22310004;
			9'd249 : dout <= 32'h1632fffd;
			9'd250 : dout <= 32'hae690000;
			9'd251 : dout <= 32'h00000000;
			9'd252 : dout <= 32'h2402000a;
			9'd253 : dout <= 32'h0000000c;
			default : dout <= 32'h0;
		endcase
	end
endmodule
